
module transkoderADC(Y,A);
input [7:0] A;
output [7:0] Y;
reg [7:0] Y;

always @(A)
case (A)
8'b00111000 : Y <=8'b00000000; // 0
8'b00111001 : Y <=8'b00000001; // 1
8'b00111010 : Y <=8'b00000010; // 2
8'b00111011 : Y <=8'b00000011; // 3
8'b00111100 : Y <=8'b00000100; // 4
8'b00111101 : Y <=8'b00000101; // 5
8'b00111110 : Y <=8'b00000110; // 6
8'b00111111 : Y <=8'b00000111; // 7
8'b01000000 : Y <=8'b00001000; // 8
8'b01000001 : Y <=8'b00001001; // 9

8'b01000010 : Y <=8'b00010000; // 10
8'b01000011 : Y <=8'b00010001; // 11
8'b01000100 : Y <=8'b00010010; // 12
8'b01000101 : Y <=8'b00010011; // 13
8'b01000110 : Y <=8'b00010100; // 14
8'b01000111 : Y <=8'b00010101; // 15
8'b01001000 : Y <=8'b00010110; // 16
8'b01001001 : Y <=8'b00010111; // 17
8'b01001010 : Y <=8'b00011000; // 18
8'b01001011 : Y <=8'b00011001; // 19

8'b01001100 : Y <=8'b00100000; // 20
8'b01001101 : Y <=8'b00100001; // 21
8'b01001110 : Y <=8'b00100010; // 22
8'b01001111 : Y <=8'b00100011; // 23
8'b01010000 : Y <=8'b00100100; // 24
8'b01010001 : Y <=8'b00100101; // 25
8'b01010010 : Y <=8'b00100110; // 26
8'b01010011 : Y <=8'b00100111; // 27
8'b01010100 : Y <=8'b00101000; // 28
8'b01010101 : Y <=8'b00101001; // 29

8'b01010110 : Y <=8'b00110000; // 30
8'b01010111 : Y <=8'b00110001; // 31
8'b01011000 : Y <=8'b00110010; // 32
8'b01011001 : Y <=8'b00110011; // 33
8'b01011010 : Y <=8'b00110100; // 34
8'b01011011 : Y <=8'b00110101; // 35
8'b01011100 : Y <=8'b00110110; // 36
8'b01011101 : Y <=8'b00110111; // 37
8'b01011110 : Y <=8'b00111000; // 38
8'b01011111 : Y <=8'b00111001; // 39

8'b01100000 : Y <=8'b01000000; // 40
8'b01100001 : Y <=8'b01000001; // 41
8'b01100010 : Y <=8'b01000010; // 42
8'b01100011 : Y <=8'b01000011; // 43
8'b01100100 : Y <=8'b01000100; // 44
8'b01100101 : Y <=8'b01000101; // 45
8'b01100110 : Y <=8'b01000110; // 46
8'b01100111 : Y <=8'b01000111; // 47
8'b01101000 : Y <=8'b01001000; // 48
8'b01101001 : Y <=8'b01001001; // 49

8'b01101010 : Y <=8'b01010000; // 50
8'b01101011 : Y <=8'b01010001; // 51
8'b01101100 : Y <=8'b01010010; // 52
8'b01101101 : Y <=8'b01010011; // 53
8'b01101110 : Y <=8'b01010100; // 54
8'b01101111 : Y <=8'b01010101; // 55
8'b01110000 : Y <=8'b01010110; // 56
8'b01110001 : Y <=8'b01010111; // 57
8'b01110010 : Y <=8'b01011000; // 58
8'b01110011 : Y <=8'b01011001; // 59

8'b01110100 : Y <=8'b01100000; // 60
8'b01110101 : Y <=8'b01100001; // 61
8'b01110110 : Y <=8'b01100010; // 62
8'b01110111 : Y <=8'b01100011; // 63
8'b01111000 : Y <=8'b01100100; // 64
8'b01111001 : Y <=8'b01100101; // 65
8'b01111010 : Y <=8'b01100110; // 66
8'b01111011 : Y <=8'b01100111; // 67
8'b01111100 : Y <=8'b01101000; // 68
8'b01111101 : Y <=8'b01101001; // 69

8'b01111110 : Y <=8'b01110000; // 70
8'b01111111 : Y <=8'b01110001; // 71
8'b10000000 : Y <=8'b01110010; // 72
8'b10000001 : Y <=8'b01110011; // 73
8'b10000010 : Y <=8'b01110100; // 74
8'b10000011 : Y <=8'b01110101; // 75
8'b10000100 : Y <=8'b01110110; // 76
8'b10000101 : Y <=8'b01110111; // 77
8'b10000110 : Y <=8'b01111000; // 78
8'b10000111 : Y <=8'b01111001; // 79

8'b10001000 : Y <=8'b10000000; // 80
8'b10001001 : Y <=8'b10000001; // 81
8'b10001010 : Y <=8'b10000010; // 82
8'b10001011 : Y <=8'b10000011; // 83
8'b10001100 : Y <=8'b10000100; // 84
8'b10001101 : Y <=8'b10000101; // 85
8'b10001110 : Y <=8'b10000110; // 86
8'b10001111 : Y <=8'b10000111; // 87
8'b10010000 : Y <=8'b10001000; // 88
8'b10010001 : Y <=8'b10001001; // 89

8'b10010010 : Y <=8'b10010000; // 90
8'b10010011 : Y <=8'b10010001; // 91
8'b10010100 : Y <=8'b10010010; // 92
8'b10010101 : Y <=8'b10010011; // 93
8'b10010110 : Y <=8'b10010100; // 94
8'b10010111 : Y <=8'b10010101; // 95
8'b10011000 : Y <=8'b10010110; // 96
8'b10011001 : Y <=8'b10010111; // 97
8'b10011010 : Y <=8'b10011000; // 98
8'b10011011 : Y <=8'b10011001; // 99
default     : Y <=8'b00100011; // 23
endcase

endmodule
