module term(WY,WE);
input [7:0] WE;
output [7:0] WY;
reg [[7:0] WY;

always @(WE)



endmodule
