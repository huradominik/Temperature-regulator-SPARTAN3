
module transkoder(Y,A);
input [7:0] A;
output [11:0] Y;
reg [11:0] Y;

always @(A)
case (A)
8'b00000000 : Y <=12'b0000_0000_0000;
8'b00000001 : Y <=12'b0000_0000_0001;
8'b00000010 : Y <=12'b0000_0000_0010;
8'b00000011 : Y <=12'b0000_0000_0011;
8'b00000100 : Y <=12'b0000_0000_0100;
8'b00000101 : Y <=12'b0000_0000_0101;
8'b00000110 : Y <=12'b0000_0000_0110;
8'b00000111 : Y <=12'b0000_0000_0111;
8'b00001000 : Y <=12'b0000_0000_1000;
8'b00001001 : Y <=12'b0000_0000_1001;

8'b00010000 : Y <=12'b0000_0001_0000;
8'b00010001 : Y <=12'b0000_0001_0001;
8'b00010010 : Y <=12'b0000_0001_0010;
8'b00010011 : Y <=12'b0000_0001_0011;
8'b00010100 : Y <=12'b0000_0001_0100;
8'b00010101 : Y <=12'b0000_0001_0101;
8'b00010110 : Y <=12'b0000_0001_0110;
8'b00010111 : Y <=12'b0000_0001_0111;
8'b00011000 : Y <=12'b0000_0001_1000;
8'b00011001 : Y <=12'b0000_0001_1001;

8'b00100000 : Y <=12'b0000_0010_0000;
8'b00100001 : Y <=12'b0000_0010_0001;
8'b00100010 : Y <=12'b0000_0010_0010;
8'b00100011 : Y <=12'b0000_0010_0011;
8'b00100100 : Y <=12'b0000_0010_0100;
8'b00100101 : Y <=12'b0000_0010_0101;
8'b00100110 : Y <=12'b0000_0010_0110;
8'b00100111 : Y <=12'b0000_0010_0111;
8'b00101000 : Y <=12'b0000_0010_1000;
8'b00101001 : Y <=12'b0000_0010_1001;

8'b00110000 : Y <=12'b0000_0011_0000;
8'b00110001 : Y <=12'b0000_0011_0001;
8'b00110010 : Y <=12'b0000_0011_0010;
8'b00110011 : Y <=12'b0000_0011_0011;
8'b00110100 : Y <=12'b0000_0011_0100;
8'b00110101 : Y <=12'b0000_0011_0101;
8'b00110110 : Y <=12'b0000_0011_0110;
8'b00110111 : Y <=12'b0000_0011_0111;
8'b00111000 : Y <=12'b0000_0011_1000;
8'b00111001 : Y <=12'b0000_0011_1001;

8'b01000000 : Y <=12'b0000_0100_0000;
8'b01000001 : Y <=12'b0000_0100_0001;
8'b01000010 : Y <=12'b0000_0100_0010;
8'b01000011 : Y <=12'b0000_0100_0011;
8'b01000100 : Y <=12'b0000_0100_0100;
8'b01000101 : Y <=12'b0000_0100_0101;
8'b01000110 : Y <=12'b0000_0100_0110;
8'b01000111 : Y <=12'b0000_0100_0111;
8'b01001000 : Y <=12'b0000_0100_1000;
8'b01001001 : Y <=12'b0000_0100_1001;

8'b01010000 : Y <=12'b0000_0101_0000;
8'b01010001 : Y <=12'b0000_0101_0001;
8'b01010010 : Y <=12'b0000_0101_0010;
8'b01010011 : Y <=12'b0000_0101_0011;
8'b01010100 : Y <=12'b0000_0101_0100;
8'b01010101 : Y <=12'b0000_0101_0101;
8'b01010110 : Y <=12'b0000_0101_0110;
8'b01010111 : Y <=12'b0000_0101_0111;
8'b01011000 : Y <=12'b0000_0101_1000;
8'b01011001 : Y <=12'b0000_0101_1001;

8'b01100000 : Y <=12'b0000_0110_0000;
8'b01100001 : Y <=12'b0000_0110_0001;
8'b01100010 : Y <=12'b0000_0110_0010;
8'b01100011 : Y <=12'b0000_0110_0011;
8'b01100100 : Y <=12'b0000_0110_0100;
8'b01100101 : Y <=12'b0000_0110_0101;
8'b01100110 : Y <=12'b0000_0110_0110;
8'b01100111 : Y <=12'b0000_0110_0111;
8'b01101000 : Y <=12'b0000_0110_1000;
8'b01101001 : Y <=12'b0000_0110_1001;

8'b01110000 : Y <=12'b0000_0111_0000;
8'b01110001 : Y <=12'b0000_0111_0001;
8'b01110010 : Y <=12'b0000_0111_0010;
8'b01110011 : Y <=12'b0000_0111_0011;
8'b01110100 : Y <=12'b0000_0111_0100;
8'b01110101 : Y <=12'b0000_0111_0101;
8'b01110110 : Y <=12'b0000_0111_0110;
8'b01110111 : Y <=12'b0000_0111_0111;
8'b01111000 : Y <=12'b0000_0111_1000;
8'b01111001 : Y <=12'b0000_0111_1001;

8'b10000000 : Y <=12'b0000_1000_0000;
8'b10000001 : Y <=12'b0000_1000_0001;
8'b10000010 : Y <=12'b0000_1000_0010;
8'b10000011 : Y <=12'b0000_1000_0011;
8'b10000100 : Y <=12'b0000_1000_0100;
8'b10000101 : Y <=12'b0000_1000_0101;
8'b10000110 : Y <=12'b0000_1000_0110;
8'b10000111 : Y <=12'b0000_1000_0111;
8'b10001000 : Y <=12'b0000_1000_1000;
8'b10001001 : Y <=12'b0000_1000_1001;

8'b10010000 : Y <=12'b0000_1001_0000;
8'b10010001 : Y <=12'b0000_1001_0001;
8'b10010010 : Y <=12'b0000_1001_0010;
8'b10010011 : Y <=12'b0000_1001_0011;
8'b10010100 : Y <=12'b0000_1001_0100;
8'b10010101 : Y <=12'b0000_1001_0101;
8'b10010110 : Y <=12'b0000_1001_0110;
8'b10010111 : Y <=12'b0000_1001_0111;
8'b10011000 : Y <=12'b0000_1001_1000;
8'b10011001 : Y <=12'b0000_1001_1001;
default : Y <=12'b0000_0011_0101;
endcase

endmodule
